
-- Autor: Marcelo Rezin
-- Data: 13/04/2020

-- Libs
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entidade
entity detector_passagem_zero is
    port(
        clock	            :   in  std_logic;
        passagem_zero       :   in  std_logic;
   
        out_display_unidade :   out std_logic_vector(6 downto 0);
        out_display_dezena  :   out std_logic_vector(6 downto 0);
        out_display_centena :   out std_logic_vector(6 downto 0);
    );
end detector_passagem_zero;

architecture main of detector_passagem_zero is

    component sete_seg_display is
        port(
            digito      :   in std_logic_vector(3 downto 0); -- valor entre 0 e 9
            out_display :   out std_logic_vector(6 downto 0)
        );
    end component sete_seg_display;

    signal unidade          :   unsigned(3 downto 0)    :=  (others => '0');
    signal dezena           :   unsigned(3 downto 0)    :=  (others => '0');
    signal centena          :   unsigned(3 downto 0)    :=  (others => '0');
    signal deteccao_zero    :   std_logic               :=  '0';
    signal reset            :   std_logic               :=  '0';

begin

    display_unidade : sete_seg_display port map (std_logic_vector(unidade), out_display_unidade);
    display_dezena  : sete_seg_display port map (std_logic_vector(dezena), out_display_dezena);
    display_centena : sete_seg_display port map (std_logic_vector(centena), out_display_centena);
	 
    process(clock)
        variable count          :   integer range 0 to 50000000 :=  0;
        variable unidade_tmp    :   unsigned(3 downto 0)    :=  (others => '0');
        variable dezena_tmp     :   unsigned(3 downto 0)    :=  (others => '0');
        variable centena_tmp    :   unsigned(3 downto 0)    :=  (others => '0');
    begin
       if rising_edge(clock) then
            count := count + 1;

            if count = 50000000 then
            --if count = 50 then
                count   :=  0; 

                unidade <=  unidade_tmp;
                dezena  <=  dezena_tmp;
                centena <=  centena_tmp;

                unidade_tmp :=  (others => '0');
                dezena_tmp  :=  (others => '0');
                centena_tmp :=  (others => '0');

                soma_tmp    <=  (others => '0');

                z   <=  '1';

            end if;

            if reset = '1' then
                reset   <=  '0';
            end if;

            if(deteccao_zero = '1') then
                reset   <=  '1';
				
                if(unidade_tmp=9) then
                    unidade_tmp :=  (others => '0');

                    if(dezena_tmp=9)then
                        dezena_tmp  :=  (others => '0');

                        centena_tmp :=  centena_tmp + 1;

                    else dezena_tmp  :=  dezena_tmp + 1;
                    end if;

                else unidade_tmp := unidade_tmp + 1;
                end if;
            end if;
       end if;

    end process;
    
    process(passagem_zero, reset)
    begin
        if reset='1' then
            deteccao_zero   <=    '0';
        elsif rising_edge(passagem_zero) then
            deteccao_zero   <=  '1';
        end if;

    end process;

end main;
